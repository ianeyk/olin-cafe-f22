`define RS2_START 24
`define RS2_END 20

`define RS1_START 19
`define RS1_END 15

`define FUNCT3_START 14
`define FUNCT3_END 12

`define FUNCT3_START 31
`define FUNCT3_END 25

`define OP_START 6
`define OP_END 0

`define RS1_START 19
`define RS1_END 15

`define RD_START 11
`define RS2_END 7

`define I_TYPE_IMM_START 31
`define I_TYPE_IMM_END 20

`define S_TYPE_IMM_1_START 31
`define S_TYPE_IMM_1_END 25

`define S_TYPE_IMM_2_START 11
`define S_TYPE_IMM_2_END 7

`define B_TYPE_IMM_1_START 31
`define B_TYPE_IMM_1_END 25

`define B_TYPE_IMM_2_START 11
`define B_TYPE_IMM_2_END 7

`define U_TYPE_IMM_START 31
`define U_TYPE_IMM_END 12

`define J_TYPE_IMM_START 31
`define J_TYPE_IMM_END 12