`ifndef INCLUDE_INSTRUCTION_DEFINES
`define INCLUDE_INSTRUCTION_DEFINES

`define RS2_START 5'd24
`define RS2_END 5'd20

`define RS1_START 5'd19
`define RS1_END 5'd15

`define FUNCT3_START 5'd14
`define FUNCT3_END 5'd12

`define FUNCT7_START 5'd31
`define FUNCT7_END 5'd25

`define OP_START 5'd6
`define OP_END 5'd0

`define RS1_START 5'd19
`define RS1_END 5'd15

`define RD_START 5'd11
`define RD_END 5'd7

`define I_TYPE_IMM_START 5'd31
`define I_TYPE_IMM_END 5'd20

`define S_TYPE_IMM_1_START 5'd31
`define S_TYPE_IMM_1_END 5'd25

`define S_TYPE_IMM_2_START 5'd11
`define S_TYPE_IMM_2_END 5'd7

`define B_TYPE_IMM_1_START 5'd31
`define B_TYPE_IMM_1_END 5'd25

`define B_TYPE_IMM_2_START 5'd11
`define B_TYPE_IMM_2_END 5'd7

`define U_TYPE_IMM_START 5'd31
`define U_TYPE_IMM_END 5'd12

`define J_TYPE_IMM_START 5'd31
`define J_TYPE_IMM_END 5'd12

`endif // INCLUDE